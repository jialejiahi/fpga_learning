/* This is a test */

module (param1, param2)
input param1;
output param2;

param2 <= param1;
endmodule
